// Computer_System.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module Computer_System (
		input  wire [8:0]   done_sram_s1_address,            //         done_sram_s1.address
		input  wire         done_sram_s1_clken,              //                     .clken
		input  wire         done_sram_s1_chipselect,         //                     .chipselect
		input  wire         done_sram_s1_write,              //                     .write
		output wire [7:0]   done_sram_s1_readdata,           //                     .readdata
		input  wire [7:0]   done_sram_s1_writedata,          //                     .writedata
		output wire         hps_io_hps_io_emac1_inst_TX_CLK, //               hps_io.hps_io_emac1_inst_TX_CLK
		output wire         hps_io_hps_io_emac1_inst_TXD0,   //                     .hps_io_emac1_inst_TXD0
		output wire         hps_io_hps_io_emac1_inst_TXD1,   //                     .hps_io_emac1_inst_TXD1
		output wire         hps_io_hps_io_emac1_inst_TXD2,   //                     .hps_io_emac1_inst_TXD2
		output wire         hps_io_hps_io_emac1_inst_TXD3,   //                     .hps_io_emac1_inst_TXD3
		input  wire         hps_io_hps_io_emac1_inst_RXD0,   //                     .hps_io_emac1_inst_RXD0
		inout  wire         hps_io_hps_io_emac1_inst_MDIO,   //                     .hps_io_emac1_inst_MDIO
		output wire         hps_io_hps_io_emac1_inst_MDC,    //                     .hps_io_emac1_inst_MDC
		input  wire         hps_io_hps_io_emac1_inst_RX_CTL, //                     .hps_io_emac1_inst_RX_CTL
		output wire         hps_io_hps_io_emac1_inst_TX_CTL, //                     .hps_io_emac1_inst_TX_CTL
		input  wire         hps_io_hps_io_emac1_inst_RX_CLK, //                     .hps_io_emac1_inst_RX_CLK
		input  wire         hps_io_hps_io_emac1_inst_RXD1,   //                     .hps_io_emac1_inst_RXD1
		input  wire         hps_io_hps_io_emac1_inst_RXD2,   //                     .hps_io_emac1_inst_RXD2
		input  wire         hps_io_hps_io_emac1_inst_RXD3,   //                     .hps_io_emac1_inst_RXD3
		inout  wire         hps_io_hps_io_qspi_inst_IO0,     //                     .hps_io_qspi_inst_IO0
		inout  wire         hps_io_hps_io_qspi_inst_IO1,     //                     .hps_io_qspi_inst_IO1
		inout  wire         hps_io_hps_io_qspi_inst_IO2,     //                     .hps_io_qspi_inst_IO2
		inout  wire         hps_io_hps_io_qspi_inst_IO3,     //                     .hps_io_qspi_inst_IO3
		output wire         hps_io_hps_io_qspi_inst_SS0,     //                     .hps_io_qspi_inst_SS0
		output wire         hps_io_hps_io_qspi_inst_CLK,     //                     .hps_io_qspi_inst_CLK
		inout  wire         hps_io_hps_io_sdio_inst_CMD,     //                     .hps_io_sdio_inst_CMD
		inout  wire         hps_io_hps_io_sdio_inst_D0,      //                     .hps_io_sdio_inst_D0
		inout  wire         hps_io_hps_io_sdio_inst_D1,      //                     .hps_io_sdio_inst_D1
		output wire         hps_io_hps_io_sdio_inst_CLK,     //                     .hps_io_sdio_inst_CLK
		inout  wire         hps_io_hps_io_sdio_inst_D2,      //                     .hps_io_sdio_inst_D2
		inout  wire         hps_io_hps_io_sdio_inst_D3,      //                     .hps_io_sdio_inst_D3
		inout  wire         hps_io_hps_io_usb1_inst_D0,      //                     .hps_io_usb1_inst_D0
		inout  wire         hps_io_hps_io_usb1_inst_D1,      //                     .hps_io_usb1_inst_D1
		inout  wire         hps_io_hps_io_usb1_inst_D2,      //                     .hps_io_usb1_inst_D2
		inout  wire         hps_io_hps_io_usb1_inst_D3,      //                     .hps_io_usb1_inst_D3
		inout  wire         hps_io_hps_io_usb1_inst_D4,      //                     .hps_io_usb1_inst_D4
		inout  wire         hps_io_hps_io_usb1_inst_D5,      //                     .hps_io_usb1_inst_D5
		inout  wire         hps_io_hps_io_usb1_inst_D6,      //                     .hps_io_usb1_inst_D6
		inout  wire         hps_io_hps_io_usb1_inst_D7,      //                     .hps_io_usb1_inst_D7
		input  wire         hps_io_hps_io_usb1_inst_CLK,     //                     .hps_io_usb1_inst_CLK
		output wire         hps_io_hps_io_usb1_inst_STP,     //                     .hps_io_usb1_inst_STP
		input  wire         hps_io_hps_io_usb1_inst_DIR,     //                     .hps_io_usb1_inst_DIR
		input  wire         hps_io_hps_io_usb1_inst_NXT,     //                     .hps_io_usb1_inst_NXT
		output wire         hps_io_hps_io_spim1_inst_CLK,    //                     .hps_io_spim1_inst_CLK
		output wire         hps_io_hps_io_spim1_inst_MOSI,   //                     .hps_io_spim1_inst_MOSI
		input  wire         hps_io_hps_io_spim1_inst_MISO,   //                     .hps_io_spim1_inst_MISO
		output wire         hps_io_hps_io_spim1_inst_SS0,    //                     .hps_io_spim1_inst_SS0
		input  wire         hps_io_hps_io_uart0_inst_RX,     //                     .hps_io_uart0_inst_RX
		output wire         hps_io_hps_io_uart0_inst_TX,     //                     .hps_io_uart0_inst_TX
		inout  wire         hps_io_hps_io_i2c0_inst_SDA,     //                     .hps_io_i2c0_inst_SDA
		inout  wire         hps_io_hps_io_i2c0_inst_SCL,     //                     .hps_io_i2c0_inst_SCL
		inout  wire         hps_io_hps_io_i2c1_inst_SDA,     //                     .hps_io_i2c1_inst_SDA
		inout  wire         hps_io_hps_io_i2c1_inst_SCL,     //                     .hps_io_i2c1_inst_SCL
		inout  wire         hps_io_hps_io_gpio_inst_GPIO09,  //                     .hps_io_gpio_inst_GPIO09
		inout  wire         hps_io_hps_io_gpio_inst_GPIO35,  //                     .hps_io_gpio_inst_GPIO35
		inout  wire         hps_io_hps_io_gpio_inst_GPIO40,  //                     .hps_io_gpio_inst_GPIO40
		inout  wire         hps_io_hps_io_gpio_inst_GPIO41,  //                     .hps_io_gpio_inst_GPIO41
		inout  wire         hps_io_hps_io_gpio_inst_GPIO48,  //                     .hps_io_gpio_inst_GPIO48
		inout  wire         hps_io_hps_io_gpio_inst_GPIO53,  //                     .hps_io_gpio_inst_GPIO53
		inout  wire         hps_io_hps_io_gpio_inst_GPIO54,  //                     .hps_io_gpio_inst_GPIO54
		inout  wire         hps_io_hps_io_gpio_inst_GPIO61,  //                     .hps_io_gpio_inst_GPIO61
		input  wire [8:0]   inst_sram_s1_address,            //         inst_sram_s1.address
		input  wire         inst_sram_s1_clken,              //                     .clken
		input  wire         inst_sram_s1_chipselect,         //                     .chipselect
		input  wire         inst_sram_s1_write,              //                     .write
		output wire [127:0] inst_sram_s1_readdata,           //                     .readdata
		input  wire [127:0] inst_sram_s1_writedata,          //                     .writedata
		input  wire [15:0]  inst_sram_s1_byteenable,         //                     .byteenable
		output wire [14:0]  memory_mem_a,                    //               memory.mem_a
		output wire [2:0]   memory_mem_ba,                   //                     .mem_ba
		output wire         memory_mem_ck,                   //                     .mem_ck
		output wire         memory_mem_ck_n,                 //                     .mem_ck_n
		output wire         memory_mem_cke,                  //                     .mem_cke
		output wire         memory_mem_cs_n,                 //                     .mem_cs_n
		output wire         memory_mem_ras_n,                //                     .mem_ras_n
		output wire         memory_mem_cas_n,                //                     .mem_cas_n
		output wire         memory_mem_we_n,                 //                     .mem_we_n
		output wire         memory_mem_reset_n,              //                     .mem_reset_n
		inout  wire [31:0]  memory_mem_dq,                   //                     .mem_dq
		inout  wire [3:0]   memory_mem_dqs,                  //                     .mem_dqs
		inout  wire [3:0]   memory_mem_dqs_n,                //                     .mem_dqs_n
		output wire         memory_mem_odt,                  //                     .mem_odt
		output wire [3:0]   memory_mem_dm,                   //                     .mem_dm
		input  wire         memory_oct_rzqin,                //                     .oct_rzqin
		input  wire         pll_0_refclk_clk,                //         pll_0_refclk.clk
		input  wire         pll_0_reset_reset,               //          pll_0_reset.reset
		output wire         sdram_clk_clk,                   //            sdram_clk.clk
		input  wire [13:0]  sram_0_s1_address,               //            sram_0_s1.address
		input  wire         sram_0_s1_clken,                 //                     .clken
		input  wire         sram_0_s1_chipselect,            //                     .chipselect
		input  wire         sram_0_s1_write,                 //                     .write
		output wire [15:0]  sram_0_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_0_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_0_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_1_s1_address,               //            sram_1_s1.address
		input  wire         sram_1_s1_clken,                 //                     .clken
		input  wire         sram_1_s1_chipselect,            //                     .chipselect
		input  wire         sram_1_s1_write,                 //                     .write
		output wire [15:0]  sram_1_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_1_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_1_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_2_s1_address,               //            sram_2_s1.address
		input  wire         sram_2_s1_clken,                 //                     .clken
		input  wire         sram_2_s1_chipselect,            //                     .chipselect
		input  wire         sram_2_s1_write,                 //                     .write
		output wire [15:0]  sram_2_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_2_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_2_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_3_s1_address,               //            sram_3_s1.address
		input  wire         sram_3_s1_clken,                 //                     .clken
		input  wire         sram_3_s1_chipselect,            //                     .chipselect
		input  wire         sram_3_s1_write,                 //                     .write
		output wire [15:0]  sram_3_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_3_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_3_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_4_s1_address,               //            sram_4_s1.address
		input  wire         sram_4_s1_clken,                 //                     .clken
		input  wire         sram_4_s1_chipselect,            //                     .chipselect
		input  wire         sram_4_s1_write,                 //                     .write
		output wire [15:0]  sram_4_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_4_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_4_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_5_s1_address,               //            sram_5_s1.address
		input  wire         sram_5_s1_clken,                 //                     .clken
		input  wire         sram_5_s1_chipselect,            //                     .chipselect
		input  wire         sram_5_s1_write,                 //                     .write
		output wire [15:0]  sram_5_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_5_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_5_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_6_s1_address,               //            sram_6_s1.address
		input  wire         sram_6_s1_clken,                 //                     .clken
		input  wire         sram_6_s1_chipselect,            //                     .chipselect
		input  wire         sram_6_s1_write,                 //                     .write
		output wire [15:0]  sram_6_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_6_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_6_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_7_s1_address,               //            sram_7_s1.address
		input  wire         sram_7_s1_clken,                 //                     .clken
		input  wire         sram_7_s1_chipselect,            //                     .chipselect
		input  wire         sram_7_s1_write,                 //                     .write
		output wire [15:0]  sram_7_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_7_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_7_s1_byteenable,            //                     .byteenable
		input  wire [13:0]  sram_8_s1_address,               //            sram_8_s1.address
		input  wire         sram_8_s1_clken,                 //                     .clken
		input  wire         sram_8_s1_chipselect,            //                     .chipselect
		input  wire         sram_8_s1_write,                 //                     .write
		output wire [15:0]  sram_8_s1_readdata,              //                     .readdata
		input  wire [15:0]  sram_8_s1_writedata,             //                     .writedata
		input  wire [1:0]   sram_8_s1_byteenable,            //                     .byteenable
		input  wire         system_pll_ref_clk_clk,          //   system_pll_ref_clk.clk
		input  wire         system_pll_ref_reset_reset       // system_pll_ref_reset.reset
	);

	wire          pll_0_outclk0_clk;                         // pll_0:outclk_0 -> [done_sram:clk, inst_sram:clk, rst_controller:clk, sram_0:clk, sram_1:clk, sram_2:clk, sram_3:clk, sram_4:clk, sram_5:clk, sram_6:clk, sram_7:clk, sram_8:clk]
	wire          system_pll_sys_clk_clk;                    // System_PLL:sys_clk_clk -> [ARM_A9_HPS:f2h_axi_clk, ARM_A9_HPS:h2f_axi_clk, ARM_A9_HPS:h2f_lw_axi_clk, done_sram:clk2, inst_sram:clk2, mm_interconnect_0:System_PLL_sys_clk_clk, rst_controller_001:clk, rst_controller_002:clk, sram_0:clk2, sram_1:clk2, sram_2:clk2, sram_3:clk2, sram_4:clk2, sram_5:clk2, sram_6:clk2, sram_7:clk2, sram_8:clk2]
	wire    [1:0] arm_a9_hps_h2f_axi_master_awburst;         // ARM_A9_HPS:h2f_AWBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awburst
	wire    [3:0] arm_a9_hps_h2f_axi_master_arlen;           // ARM_A9_HPS:h2f_ARLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlen
	wire   [15:0] arm_a9_hps_h2f_axi_master_wstrb;           // ARM_A9_HPS:h2f_WSTRB -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wstrb
	wire          arm_a9_hps_h2f_axi_master_wready;          // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wready -> ARM_A9_HPS:h2f_WREADY
	wire   [11:0] arm_a9_hps_h2f_axi_master_rid;             // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rid -> ARM_A9_HPS:h2f_RID
	wire          arm_a9_hps_h2f_axi_master_rready;          // ARM_A9_HPS:h2f_RREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rready
	wire    [3:0] arm_a9_hps_h2f_axi_master_awlen;           // ARM_A9_HPS:h2f_AWLEN -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlen
	wire   [11:0] arm_a9_hps_h2f_axi_master_wid;             // ARM_A9_HPS:h2f_WID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wid
	wire    [3:0] arm_a9_hps_h2f_axi_master_arcache;         // ARM_A9_HPS:h2f_ARCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arcache
	wire          arm_a9_hps_h2f_axi_master_wvalid;          // ARM_A9_HPS:h2f_WVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wvalid
	wire   [29:0] arm_a9_hps_h2f_axi_master_araddr;          // ARM_A9_HPS:h2f_ARADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_araddr
	wire    [2:0] arm_a9_hps_h2f_axi_master_arprot;          // ARM_A9_HPS:h2f_ARPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arprot
	wire    [2:0] arm_a9_hps_h2f_axi_master_awprot;          // ARM_A9_HPS:h2f_AWPROT -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awprot
	wire  [127:0] arm_a9_hps_h2f_axi_master_wdata;           // ARM_A9_HPS:h2f_WDATA -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wdata
	wire          arm_a9_hps_h2f_axi_master_arvalid;         // ARM_A9_HPS:h2f_ARVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arvalid
	wire    [3:0] arm_a9_hps_h2f_axi_master_awcache;         // ARM_A9_HPS:h2f_AWCACHE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awcache
	wire   [11:0] arm_a9_hps_h2f_axi_master_arid;            // ARM_A9_HPS:h2f_ARID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arid
	wire    [1:0] arm_a9_hps_h2f_axi_master_arlock;          // ARM_A9_HPS:h2f_ARLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arlock
	wire    [1:0] arm_a9_hps_h2f_axi_master_awlock;          // ARM_A9_HPS:h2f_AWLOCK -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awlock
	wire   [29:0] arm_a9_hps_h2f_axi_master_awaddr;          // ARM_A9_HPS:h2f_AWADDR -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awaddr
	wire    [1:0] arm_a9_hps_h2f_axi_master_bresp;           // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bresp -> ARM_A9_HPS:h2f_BRESP
	wire          arm_a9_hps_h2f_axi_master_arready;         // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arready -> ARM_A9_HPS:h2f_ARREADY
	wire  [127:0] arm_a9_hps_h2f_axi_master_rdata;           // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rdata -> ARM_A9_HPS:h2f_RDATA
	wire          arm_a9_hps_h2f_axi_master_awready;         // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awready -> ARM_A9_HPS:h2f_AWREADY
	wire    [1:0] arm_a9_hps_h2f_axi_master_arburst;         // ARM_A9_HPS:h2f_ARBURST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arburst
	wire    [2:0] arm_a9_hps_h2f_axi_master_arsize;          // ARM_A9_HPS:h2f_ARSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_arsize
	wire          arm_a9_hps_h2f_axi_master_bready;          // ARM_A9_HPS:h2f_BREADY -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bready
	wire          arm_a9_hps_h2f_axi_master_rlast;           // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rlast -> ARM_A9_HPS:h2f_RLAST
	wire          arm_a9_hps_h2f_axi_master_wlast;           // ARM_A9_HPS:h2f_WLAST -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_wlast
	wire    [1:0] arm_a9_hps_h2f_axi_master_rresp;           // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rresp -> ARM_A9_HPS:h2f_RRESP
	wire   [11:0] arm_a9_hps_h2f_axi_master_awid;            // ARM_A9_HPS:h2f_AWID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awid
	wire   [11:0] arm_a9_hps_h2f_axi_master_bid;             // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bid -> ARM_A9_HPS:h2f_BID
	wire          arm_a9_hps_h2f_axi_master_bvalid;          // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_bvalid -> ARM_A9_HPS:h2f_BVALID
	wire    [2:0] arm_a9_hps_h2f_axi_master_awsize;          // ARM_A9_HPS:h2f_AWSIZE -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awsize
	wire          arm_a9_hps_h2f_axi_master_awvalid;         // ARM_A9_HPS:h2f_AWVALID -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_awvalid
	wire          arm_a9_hps_h2f_axi_master_rvalid;          // mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_rvalid -> ARM_A9_HPS:h2f_RVALID
	wire          mm_interconnect_0_inst_sram_s2_chipselect; // mm_interconnect_0:inst_sram_s2_chipselect -> inst_sram:chipselect2
	wire  [127:0] mm_interconnect_0_inst_sram_s2_readdata;   // inst_sram:readdata2 -> mm_interconnect_0:inst_sram_s2_readdata
	wire    [8:0] mm_interconnect_0_inst_sram_s2_address;    // mm_interconnect_0:inst_sram_s2_address -> inst_sram:address2
	wire   [15:0] mm_interconnect_0_inst_sram_s2_byteenable; // mm_interconnect_0:inst_sram_s2_byteenable -> inst_sram:byteenable2
	wire          mm_interconnect_0_inst_sram_s2_write;      // mm_interconnect_0:inst_sram_s2_write -> inst_sram:write2
	wire  [127:0] mm_interconnect_0_inst_sram_s2_writedata;  // mm_interconnect_0:inst_sram_s2_writedata -> inst_sram:writedata2
	wire          mm_interconnect_0_inst_sram_s2_clken;      // mm_interconnect_0:inst_sram_s2_clken -> inst_sram:clken2
	wire          mm_interconnect_0_sram_0_s2_chipselect;    // mm_interconnect_0:sram_0_s2_chipselect -> sram_0:chipselect2
	wire   [15:0] mm_interconnect_0_sram_0_s2_readdata;      // sram_0:readdata2 -> mm_interconnect_0:sram_0_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_0_s2_address;       // mm_interconnect_0:sram_0_s2_address -> sram_0:address2
	wire    [1:0] mm_interconnect_0_sram_0_s2_byteenable;    // mm_interconnect_0:sram_0_s2_byteenable -> sram_0:byteenable2
	wire          mm_interconnect_0_sram_0_s2_write;         // mm_interconnect_0:sram_0_s2_write -> sram_0:write2
	wire   [15:0] mm_interconnect_0_sram_0_s2_writedata;     // mm_interconnect_0:sram_0_s2_writedata -> sram_0:writedata2
	wire          mm_interconnect_0_sram_0_s2_clken;         // mm_interconnect_0:sram_0_s2_clken -> sram_0:clken2
	wire          mm_interconnect_0_sram_1_s2_chipselect;    // mm_interconnect_0:sram_1_s2_chipselect -> sram_1:chipselect2
	wire   [15:0] mm_interconnect_0_sram_1_s2_readdata;      // sram_1:readdata2 -> mm_interconnect_0:sram_1_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_1_s2_address;       // mm_interconnect_0:sram_1_s2_address -> sram_1:address2
	wire    [1:0] mm_interconnect_0_sram_1_s2_byteenable;    // mm_interconnect_0:sram_1_s2_byteenable -> sram_1:byteenable2
	wire          mm_interconnect_0_sram_1_s2_write;         // mm_interconnect_0:sram_1_s2_write -> sram_1:write2
	wire   [15:0] mm_interconnect_0_sram_1_s2_writedata;     // mm_interconnect_0:sram_1_s2_writedata -> sram_1:writedata2
	wire          mm_interconnect_0_sram_1_s2_clken;         // mm_interconnect_0:sram_1_s2_clken -> sram_1:clken2
	wire          mm_interconnect_0_sram_2_s2_chipselect;    // mm_interconnect_0:sram_2_s2_chipselect -> sram_2:chipselect2
	wire   [15:0] mm_interconnect_0_sram_2_s2_readdata;      // sram_2:readdata2 -> mm_interconnect_0:sram_2_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_2_s2_address;       // mm_interconnect_0:sram_2_s2_address -> sram_2:address2
	wire    [1:0] mm_interconnect_0_sram_2_s2_byteenable;    // mm_interconnect_0:sram_2_s2_byteenable -> sram_2:byteenable2
	wire          mm_interconnect_0_sram_2_s2_write;         // mm_interconnect_0:sram_2_s2_write -> sram_2:write2
	wire   [15:0] mm_interconnect_0_sram_2_s2_writedata;     // mm_interconnect_0:sram_2_s2_writedata -> sram_2:writedata2
	wire          mm_interconnect_0_sram_2_s2_clken;         // mm_interconnect_0:sram_2_s2_clken -> sram_2:clken2
	wire          mm_interconnect_0_sram_3_s2_chipselect;    // mm_interconnect_0:sram_3_s2_chipselect -> sram_3:chipselect2
	wire   [15:0] mm_interconnect_0_sram_3_s2_readdata;      // sram_3:readdata2 -> mm_interconnect_0:sram_3_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_3_s2_address;       // mm_interconnect_0:sram_3_s2_address -> sram_3:address2
	wire    [1:0] mm_interconnect_0_sram_3_s2_byteenable;    // mm_interconnect_0:sram_3_s2_byteenable -> sram_3:byteenable2
	wire          mm_interconnect_0_sram_3_s2_write;         // mm_interconnect_0:sram_3_s2_write -> sram_3:write2
	wire   [15:0] mm_interconnect_0_sram_3_s2_writedata;     // mm_interconnect_0:sram_3_s2_writedata -> sram_3:writedata2
	wire          mm_interconnect_0_sram_3_s2_clken;         // mm_interconnect_0:sram_3_s2_clken -> sram_3:clken2
	wire          mm_interconnect_0_sram_4_s2_chipselect;    // mm_interconnect_0:sram_4_s2_chipselect -> sram_4:chipselect2
	wire   [15:0] mm_interconnect_0_sram_4_s2_readdata;      // sram_4:readdata2 -> mm_interconnect_0:sram_4_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_4_s2_address;       // mm_interconnect_0:sram_4_s2_address -> sram_4:address2
	wire    [1:0] mm_interconnect_0_sram_4_s2_byteenable;    // mm_interconnect_0:sram_4_s2_byteenable -> sram_4:byteenable2
	wire          mm_interconnect_0_sram_4_s2_write;         // mm_interconnect_0:sram_4_s2_write -> sram_4:write2
	wire   [15:0] mm_interconnect_0_sram_4_s2_writedata;     // mm_interconnect_0:sram_4_s2_writedata -> sram_4:writedata2
	wire          mm_interconnect_0_sram_4_s2_clken;         // mm_interconnect_0:sram_4_s2_clken -> sram_4:clken2
	wire          mm_interconnect_0_sram_5_s2_chipselect;    // mm_interconnect_0:sram_5_s2_chipselect -> sram_5:chipselect2
	wire   [15:0] mm_interconnect_0_sram_5_s2_readdata;      // sram_5:readdata2 -> mm_interconnect_0:sram_5_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_5_s2_address;       // mm_interconnect_0:sram_5_s2_address -> sram_5:address2
	wire    [1:0] mm_interconnect_0_sram_5_s2_byteenable;    // mm_interconnect_0:sram_5_s2_byteenable -> sram_5:byteenable2
	wire          mm_interconnect_0_sram_5_s2_write;         // mm_interconnect_0:sram_5_s2_write -> sram_5:write2
	wire   [15:0] mm_interconnect_0_sram_5_s2_writedata;     // mm_interconnect_0:sram_5_s2_writedata -> sram_5:writedata2
	wire          mm_interconnect_0_sram_5_s2_clken;         // mm_interconnect_0:sram_5_s2_clken -> sram_5:clken2
	wire          mm_interconnect_0_sram_6_s2_chipselect;    // mm_interconnect_0:sram_6_s2_chipselect -> sram_6:chipselect2
	wire   [15:0] mm_interconnect_0_sram_6_s2_readdata;      // sram_6:readdata2 -> mm_interconnect_0:sram_6_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_6_s2_address;       // mm_interconnect_0:sram_6_s2_address -> sram_6:address2
	wire    [1:0] mm_interconnect_0_sram_6_s2_byteenable;    // mm_interconnect_0:sram_6_s2_byteenable -> sram_6:byteenable2
	wire          mm_interconnect_0_sram_6_s2_write;         // mm_interconnect_0:sram_6_s2_write -> sram_6:write2
	wire   [15:0] mm_interconnect_0_sram_6_s2_writedata;     // mm_interconnect_0:sram_6_s2_writedata -> sram_6:writedata2
	wire          mm_interconnect_0_sram_6_s2_clken;         // mm_interconnect_0:sram_6_s2_clken -> sram_6:clken2
	wire          mm_interconnect_0_sram_7_s2_chipselect;    // mm_interconnect_0:sram_7_s2_chipselect -> sram_7:chipselect2
	wire   [15:0] mm_interconnect_0_sram_7_s2_readdata;      // sram_7:readdata2 -> mm_interconnect_0:sram_7_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_7_s2_address;       // mm_interconnect_0:sram_7_s2_address -> sram_7:address2
	wire    [1:0] mm_interconnect_0_sram_7_s2_byteenable;    // mm_interconnect_0:sram_7_s2_byteenable -> sram_7:byteenable2
	wire          mm_interconnect_0_sram_7_s2_write;         // mm_interconnect_0:sram_7_s2_write -> sram_7:write2
	wire   [15:0] mm_interconnect_0_sram_7_s2_writedata;     // mm_interconnect_0:sram_7_s2_writedata -> sram_7:writedata2
	wire          mm_interconnect_0_sram_7_s2_clken;         // mm_interconnect_0:sram_7_s2_clken -> sram_7:clken2
	wire          mm_interconnect_0_sram_8_s2_chipselect;    // mm_interconnect_0:sram_8_s2_chipselect -> sram_8:chipselect2
	wire   [15:0] mm_interconnect_0_sram_8_s2_readdata;      // sram_8:readdata2 -> mm_interconnect_0:sram_8_s2_readdata
	wire   [13:0] mm_interconnect_0_sram_8_s2_address;       // mm_interconnect_0:sram_8_s2_address -> sram_8:address2
	wire    [1:0] mm_interconnect_0_sram_8_s2_byteenable;    // mm_interconnect_0:sram_8_s2_byteenable -> sram_8:byteenable2
	wire          mm_interconnect_0_sram_8_s2_write;         // mm_interconnect_0:sram_8_s2_write -> sram_8:write2
	wire   [15:0] mm_interconnect_0_sram_8_s2_writedata;     // mm_interconnect_0:sram_8_s2_writedata -> sram_8:writedata2
	wire          mm_interconnect_0_sram_8_s2_clken;         // mm_interconnect_0:sram_8_s2_clken -> sram_8:clken2
	wire          mm_interconnect_0_done_sram_s2_chipselect; // mm_interconnect_0:done_sram_s2_chipselect -> done_sram:chipselect2
	wire    [7:0] mm_interconnect_0_done_sram_s2_readdata;   // done_sram:readdata2 -> mm_interconnect_0:done_sram_s2_readdata
	wire    [8:0] mm_interconnect_0_done_sram_s2_address;    // mm_interconnect_0:done_sram_s2_address -> done_sram:address2
	wire          mm_interconnect_0_done_sram_s2_write;      // mm_interconnect_0:done_sram_s2_write -> done_sram:write2
	wire    [7:0] mm_interconnect_0_done_sram_s2_writedata;  // mm_interconnect_0:done_sram_s2_writedata -> done_sram:writedata2
	wire          mm_interconnect_0_done_sram_s2_clken;      // mm_interconnect_0:done_sram_s2_clken -> done_sram:clken2
	wire   [31:0] arm_a9_hps_f2h_irq0_irq;                   // irq_mapper:sender_irq -> ARM_A9_HPS:f2h_irq_p0
	wire   [31:0] arm_a9_hps_f2h_irq1_irq;                   // irq_mapper_001:sender_irq -> ARM_A9_HPS:f2h_irq_p1
	wire          rst_controller_reset_out_reset;            // rst_controller:reset_out -> [done_sram:reset, inst_sram:reset, sram_0:reset, sram_1:reset, sram_2:reset, sram_3:reset, sram_4:reset, sram_5:reset, sram_6:reset, sram_7:reset, sram_8:reset]
	wire          rst_controller_reset_out_reset_req;        // rst_controller:reset_req -> [done_sram:reset_req, inst_sram:reset_req, sram_0:reset_req, sram_1:reset_req, sram_2:reset_req, sram_3:reset_req, sram_4:reset_req, sram_5:reset_req, sram_6:reset_req, sram_7:reset_req, sram_8:reset_req]
	wire          arm_a9_hps_h2f_reset_reset;                // ARM_A9_HPS:h2f_rst_n -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0]
	wire          system_pll_reset_source_reset;             // System_PLL:reset_source_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire          rst_controller_001_reset_out_reset;        // rst_controller_001:reset_out -> [done_sram:reset2, inst_sram:reset2, mm_interconnect_0:inst_sram_reset2_reset_bridge_in_reset_reset, sram_0:reset2, sram_1:reset2, sram_2:reset2, sram_3:reset2, sram_4:reset2, sram_5:reset2, sram_6:reset2, sram_7:reset2, sram_8:reset2]
	wire          rst_controller_001_reset_out_reset_req;    // rst_controller_001:reset_req -> [done_sram:reset_req2, inst_sram:reset_req2, sram_0:reset_req2, sram_1:reset_req2, sram_2:reset_req2, sram_3:reset_req2, sram_4:reset_req2, sram_5:reset_req2, sram_6:reset_req2, sram_7:reset_req2, sram_8:reset_req2]
	wire          rst_controller_002_reset_out_reset;        // rst_controller_002:reset_out -> mm_interconnect_0:ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset

	Computer_System_ARM_A9_HPS #(
		.F2S_Width (2),
		.S2F_Width (3)
	) arm_a9_hps (
		.mem_a                    (memory_mem_a),                      //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                     //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                     //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                   //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                    //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                   //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                  //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                  //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                   //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                     //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                    //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                  //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                    //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                     //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                  //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),   //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),     //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),     //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),     //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),     //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),     //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),     //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),      //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),   //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),   //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),   //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),     //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),     //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),     //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),       //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),       //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),       //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),       //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),       //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),       //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),       //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),        //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),        //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),       //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),        //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),        //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),        //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),        //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),        //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),        //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),        //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),        //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),        //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),        //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),       //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),       //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),       //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),       //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_io_hps_io_spim1_inst_CLK),      //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_io_hps_io_spim1_inst_MOSI),     //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_io_hps_io_spim1_inst_MISO),     //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_io_hps_io_spim1_inst_SS0),      //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),       //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),       //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),       //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),       //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),       //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),       //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),    //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_io_hps_io_gpio_inst_GPIO35),    //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),    //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),    //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),    //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_io_hps_io_gpio_inst_GPIO53),    //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_io_hps_io_gpio_inst_GPIO54),    //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_io_hps_io_gpio_inst_GPIO61),    //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (arm_a9_hps_h2f_reset_reset),        //         h2f_reset.reset_n
		.h2f_axi_clk              (system_pll_sys_clk_clk),            //     h2f_axi_clock.clk
		.h2f_AWID                 (arm_a9_hps_h2f_axi_master_awid),    //    h2f_axi_master.awid
		.h2f_AWADDR               (arm_a9_hps_h2f_axi_master_awaddr),  //                  .awaddr
		.h2f_AWLEN                (arm_a9_hps_h2f_axi_master_awlen),   //                  .awlen
		.h2f_AWSIZE               (arm_a9_hps_h2f_axi_master_awsize),  //                  .awsize
		.h2f_AWBURST              (arm_a9_hps_h2f_axi_master_awburst), //                  .awburst
		.h2f_AWLOCK               (arm_a9_hps_h2f_axi_master_awlock),  //                  .awlock
		.h2f_AWCACHE              (arm_a9_hps_h2f_axi_master_awcache), //                  .awcache
		.h2f_AWPROT               (arm_a9_hps_h2f_axi_master_awprot),  //                  .awprot
		.h2f_AWVALID              (arm_a9_hps_h2f_axi_master_awvalid), //                  .awvalid
		.h2f_AWREADY              (arm_a9_hps_h2f_axi_master_awready), //                  .awready
		.h2f_WID                  (arm_a9_hps_h2f_axi_master_wid),     //                  .wid
		.h2f_WDATA                (arm_a9_hps_h2f_axi_master_wdata),   //                  .wdata
		.h2f_WSTRB                (arm_a9_hps_h2f_axi_master_wstrb),   //                  .wstrb
		.h2f_WLAST                (arm_a9_hps_h2f_axi_master_wlast),   //                  .wlast
		.h2f_WVALID               (arm_a9_hps_h2f_axi_master_wvalid),  //                  .wvalid
		.h2f_WREADY               (arm_a9_hps_h2f_axi_master_wready),  //                  .wready
		.h2f_BID                  (arm_a9_hps_h2f_axi_master_bid),     //                  .bid
		.h2f_BRESP                (arm_a9_hps_h2f_axi_master_bresp),   //                  .bresp
		.h2f_BVALID               (arm_a9_hps_h2f_axi_master_bvalid),  //                  .bvalid
		.h2f_BREADY               (arm_a9_hps_h2f_axi_master_bready),  //                  .bready
		.h2f_ARID                 (arm_a9_hps_h2f_axi_master_arid),    //                  .arid
		.h2f_ARADDR               (arm_a9_hps_h2f_axi_master_araddr),  //                  .araddr
		.h2f_ARLEN                (arm_a9_hps_h2f_axi_master_arlen),   //                  .arlen
		.h2f_ARSIZE               (arm_a9_hps_h2f_axi_master_arsize),  //                  .arsize
		.h2f_ARBURST              (arm_a9_hps_h2f_axi_master_arburst), //                  .arburst
		.h2f_ARLOCK               (arm_a9_hps_h2f_axi_master_arlock),  //                  .arlock
		.h2f_ARCACHE              (arm_a9_hps_h2f_axi_master_arcache), //                  .arcache
		.h2f_ARPROT               (arm_a9_hps_h2f_axi_master_arprot),  //                  .arprot
		.h2f_ARVALID              (arm_a9_hps_h2f_axi_master_arvalid), //                  .arvalid
		.h2f_ARREADY              (arm_a9_hps_h2f_axi_master_arready), //                  .arready
		.h2f_RID                  (arm_a9_hps_h2f_axi_master_rid),     //                  .rid
		.h2f_RDATA                (arm_a9_hps_h2f_axi_master_rdata),   //                  .rdata
		.h2f_RRESP                (arm_a9_hps_h2f_axi_master_rresp),   //                  .rresp
		.h2f_RLAST                (arm_a9_hps_h2f_axi_master_rlast),   //                  .rlast
		.h2f_RVALID               (arm_a9_hps_h2f_axi_master_rvalid),  //                  .rvalid
		.h2f_RREADY               (arm_a9_hps_h2f_axi_master_rready),  //                  .rready
		.f2h_axi_clk              (system_pll_sys_clk_clk),            //     f2h_axi_clock.clk
		.f2h_AWID                 (),                                  //     f2h_axi_slave.awid
		.f2h_AWADDR               (),                                  //                  .awaddr
		.f2h_AWLEN                (),                                  //                  .awlen
		.f2h_AWSIZE               (),                                  //                  .awsize
		.f2h_AWBURST              (),                                  //                  .awburst
		.f2h_AWLOCK               (),                                  //                  .awlock
		.f2h_AWCACHE              (),                                  //                  .awcache
		.f2h_AWPROT               (),                                  //                  .awprot
		.f2h_AWVALID              (),                                  //                  .awvalid
		.f2h_AWREADY              (),                                  //                  .awready
		.f2h_AWUSER               (),                                  //                  .awuser
		.f2h_WID                  (),                                  //                  .wid
		.f2h_WDATA                (),                                  //                  .wdata
		.f2h_WSTRB                (),                                  //                  .wstrb
		.f2h_WLAST                (),                                  //                  .wlast
		.f2h_WVALID               (),                                  //                  .wvalid
		.f2h_WREADY               (),                                  //                  .wready
		.f2h_BID                  (),                                  //                  .bid
		.f2h_BRESP                (),                                  //                  .bresp
		.f2h_BVALID               (),                                  //                  .bvalid
		.f2h_BREADY               (),                                  //                  .bready
		.f2h_ARID                 (),                                  //                  .arid
		.f2h_ARADDR               (),                                  //                  .araddr
		.f2h_ARLEN                (),                                  //                  .arlen
		.f2h_ARSIZE               (),                                  //                  .arsize
		.f2h_ARBURST              (),                                  //                  .arburst
		.f2h_ARLOCK               (),                                  //                  .arlock
		.f2h_ARCACHE              (),                                  //                  .arcache
		.f2h_ARPROT               (),                                  //                  .arprot
		.f2h_ARVALID              (),                                  //                  .arvalid
		.f2h_ARREADY              (),                                  //                  .arready
		.f2h_ARUSER               (),                                  //                  .aruser
		.f2h_RID                  (),                                  //                  .rid
		.f2h_RDATA                (),                                  //                  .rdata
		.f2h_RRESP                (),                                  //                  .rresp
		.f2h_RLAST                (),                                  //                  .rlast
		.f2h_RVALID               (),                                  //                  .rvalid
		.f2h_RREADY               (),                                  //                  .rready
		.h2f_lw_axi_clk           (system_pll_sys_clk_clk),            //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (),                                  // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (),                                  //                  .awaddr
		.h2f_lw_AWLEN             (),                                  //                  .awlen
		.h2f_lw_AWSIZE            (),                                  //                  .awsize
		.h2f_lw_AWBURST           (),                                  //                  .awburst
		.h2f_lw_AWLOCK            (),                                  //                  .awlock
		.h2f_lw_AWCACHE           (),                                  //                  .awcache
		.h2f_lw_AWPROT            (),                                  //                  .awprot
		.h2f_lw_AWVALID           (),                                  //                  .awvalid
		.h2f_lw_AWREADY           (),                                  //                  .awready
		.h2f_lw_WID               (),                                  //                  .wid
		.h2f_lw_WDATA             (),                                  //                  .wdata
		.h2f_lw_WSTRB             (),                                  //                  .wstrb
		.h2f_lw_WLAST             (),                                  //                  .wlast
		.h2f_lw_WVALID            (),                                  //                  .wvalid
		.h2f_lw_WREADY            (),                                  //                  .wready
		.h2f_lw_BID               (),                                  //                  .bid
		.h2f_lw_BRESP             (),                                  //                  .bresp
		.h2f_lw_BVALID            (),                                  //                  .bvalid
		.h2f_lw_BREADY            (),                                  //                  .bready
		.h2f_lw_ARID              (),                                  //                  .arid
		.h2f_lw_ARADDR            (),                                  //                  .araddr
		.h2f_lw_ARLEN             (),                                  //                  .arlen
		.h2f_lw_ARSIZE            (),                                  //                  .arsize
		.h2f_lw_ARBURST           (),                                  //                  .arburst
		.h2f_lw_ARLOCK            (),                                  //                  .arlock
		.h2f_lw_ARCACHE           (),                                  //                  .arcache
		.h2f_lw_ARPROT            (),                                  //                  .arprot
		.h2f_lw_ARVALID           (),                                  //                  .arvalid
		.h2f_lw_ARREADY           (),                                  //                  .arready
		.h2f_lw_RID               (),                                  //                  .rid
		.h2f_lw_RDATA             (),                                  //                  .rdata
		.h2f_lw_RRESP             (),                                  //                  .rresp
		.h2f_lw_RLAST             (),                                  //                  .rlast
		.h2f_lw_RVALID            (),                                  //                  .rvalid
		.h2f_lw_RREADY            (),                                  //                  .rready
		.f2h_irq_p0               (arm_a9_hps_f2h_irq0_irq),           //          f2h_irq0.irq
		.f2h_irq_p1               (arm_a9_hps_f2h_irq1_irq)            //          f2h_irq1.irq
	);

	Computer_System_System_PLL system_pll (
		.ref_clk_clk        (system_pll_ref_clk_clk),        //      ref_clk.clk
		.ref_reset_reset    (system_pll_ref_reset_reset),    //    ref_reset.reset
		.sys_clk_clk        (system_pll_sys_clk_clk),        //      sys_clk.clk
		.sdram_clk_clk      (sdram_clk_clk),                 //    sdram_clk.clk
		.reset_source_reset (system_pll_reset_source_reset)  // reset_source.reset
	);

	Computer_System_done_sram done_sram (
		.clk         (pll_0_outclk0_clk),                         //   clk1.clk
		.address     (done_sram_s1_address),                      //     s1.address
		.clken       (done_sram_s1_clken),                        //       .clken
		.chipselect  (done_sram_s1_chipselect),                   //       .chipselect
		.write       (done_sram_s1_write),                        //       .write
		.readdata    (done_sram_s1_readdata),                     //       .readdata
		.writedata   (done_sram_s1_writedata),                    //       .writedata
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.address2    (mm_interconnect_0_done_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_done_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_done_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_done_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_done_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_done_sram_s2_writedata),  //       .writedata
		.clk2        (system_pll_sys_clk_clk),                    //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),        // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	Computer_System_inst_sram inst_sram (
		.clk         (pll_0_outclk0_clk),                         //   clk1.clk
		.address     (inst_sram_s1_address),                      //     s1.address
		.clken       (inst_sram_s1_clken),                        //       .clken
		.chipselect  (inst_sram_s1_chipselect),                   //       .chipselect
		.write       (inst_sram_s1_write),                        //       .write
		.readdata    (inst_sram_s1_readdata),                     //       .readdata
		.writedata   (inst_sram_s1_writedata),                    //       .writedata
		.byteenable  (inst_sram_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),            // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),        //       .reset_req
		.address2    (mm_interconnect_0_inst_sram_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_inst_sram_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_inst_sram_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_inst_sram_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_inst_sram_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_inst_sram_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_inst_sram_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                    //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),        // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),    //       .reset_req
		.freeze      (1'b0)                                       // (terminated)
	);

	Computer_System_pll_0 pll_0 (
		.refclk   (pll_0_refclk_clk),  //  refclk.clk
		.rst      (pll_0_reset_reset), //   reset.reset
		.outclk_0 (pll_0_outclk0_clk), // outclk0.clk
		.locked   ()                   // (terminated)
	);

	Computer_System_sram_0 sram_0 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_0_s1_address),                      //     s1.address
		.clken       (sram_0_s1_clken),                        //       .clken
		.chipselect  (sram_0_s1_chipselect),                   //       .chipselect
		.write       (sram_0_s1_write),                        //       .write
		.readdata    (sram_0_s1_readdata),                     //       .readdata
		.writedata   (sram_0_s1_writedata),                    //       .writedata
		.byteenable  (sram_0_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_0_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_0_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_0_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_0_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_0_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_0_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_0_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_1 sram_1 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_1_s1_address),                      //     s1.address
		.clken       (sram_1_s1_clken),                        //       .clken
		.chipselect  (sram_1_s1_chipselect),                   //       .chipselect
		.write       (sram_1_s1_write),                        //       .write
		.readdata    (sram_1_s1_readdata),                     //       .readdata
		.writedata   (sram_1_s1_writedata),                    //       .writedata
		.byteenable  (sram_1_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_1_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_1_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_1_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_1_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_1_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_1_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_1_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_2 sram_2 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_2_s1_address),                      //     s1.address
		.clken       (sram_2_s1_clken),                        //       .clken
		.chipselect  (sram_2_s1_chipselect),                   //       .chipselect
		.write       (sram_2_s1_write),                        //       .write
		.readdata    (sram_2_s1_readdata),                     //       .readdata
		.writedata   (sram_2_s1_writedata),                    //       .writedata
		.byteenable  (sram_2_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_2_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_2_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_2_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_2_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_2_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_2_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_2_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_3 sram_3 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_3_s1_address),                      //     s1.address
		.clken       (sram_3_s1_clken),                        //       .clken
		.chipselect  (sram_3_s1_chipselect),                   //       .chipselect
		.write       (sram_3_s1_write),                        //       .write
		.readdata    (sram_3_s1_readdata),                     //       .readdata
		.writedata   (sram_3_s1_writedata),                    //       .writedata
		.byteenable  (sram_3_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_3_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_3_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_3_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_3_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_3_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_3_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_3_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_4 sram_4 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_4_s1_address),                      //     s1.address
		.clken       (sram_4_s1_clken),                        //       .clken
		.chipselect  (sram_4_s1_chipselect),                   //       .chipselect
		.write       (sram_4_s1_write),                        //       .write
		.readdata    (sram_4_s1_readdata),                     //       .readdata
		.writedata   (sram_4_s1_writedata),                    //       .writedata
		.byteenable  (sram_4_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_4_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_4_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_4_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_4_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_4_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_4_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_4_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_5 sram_5 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_5_s1_address),                      //     s1.address
		.clken       (sram_5_s1_clken),                        //       .clken
		.chipselect  (sram_5_s1_chipselect),                   //       .chipselect
		.write       (sram_5_s1_write),                        //       .write
		.readdata    (sram_5_s1_readdata),                     //       .readdata
		.writedata   (sram_5_s1_writedata),                    //       .writedata
		.byteenable  (sram_5_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_5_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_5_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_5_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_5_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_5_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_5_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_5_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_6 sram_6 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_6_s1_address),                      //     s1.address
		.clken       (sram_6_s1_clken),                        //       .clken
		.chipselect  (sram_6_s1_chipselect),                   //       .chipselect
		.write       (sram_6_s1_write),                        //       .write
		.readdata    (sram_6_s1_readdata),                     //       .readdata
		.writedata   (sram_6_s1_writedata),                    //       .writedata
		.byteenable  (sram_6_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_6_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_6_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_6_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_6_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_6_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_6_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_6_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_7 sram_7 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_7_s1_address),                      //     s1.address
		.clken       (sram_7_s1_clken),                        //       .clken
		.chipselect  (sram_7_s1_chipselect),                   //       .chipselect
		.write       (sram_7_s1_write),                        //       .write
		.readdata    (sram_7_s1_readdata),                     //       .readdata
		.writedata   (sram_7_s1_writedata),                    //       .writedata
		.byteenable  (sram_7_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_7_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_7_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_7_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_7_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_7_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_7_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_7_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_sram_8 sram_8 (
		.clk         (pll_0_outclk0_clk),                      //   clk1.clk
		.address     (sram_8_s1_address),                      //     s1.address
		.clken       (sram_8_s1_clken),                        //       .clken
		.chipselect  (sram_8_s1_chipselect),                   //       .chipselect
		.write       (sram_8_s1_write),                        //       .write
		.readdata    (sram_8_s1_readdata),                     //       .readdata
		.writedata   (sram_8_s1_writedata),                    //       .writedata
		.byteenable  (sram_8_s1_byteenable),                   //       .byteenable
		.reset       (rst_controller_reset_out_reset),         // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),     //       .reset_req
		.address2    (mm_interconnect_0_sram_8_s2_address),    //     s2.address
		.chipselect2 (mm_interconnect_0_sram_8_s2_chipselect), //       .chipselect
		.clken2      (mm_interconnect_0_sram_8_s2_clken),      //       .clken
		.write2      (mm_interconnect_0_sram_8_s2_write),      //       .write
		.readdata2   (mm_interconnect_0_sram_8_s2_readdata),   //       .readdata
		.writedata2  (mm_interconnect_0_sram_8_s2_writedata),  //       .writedata
		.byteenable2 (mm_interconnect_0_sram_8_s2_byteenable), //       .byteenable
		.clk2        (system_pll_sys_clk_clk),                 //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),     // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze      (1'b0)                                    // (terminated)
	);

	Computer_System_mm_interconnect_0 mm_interconnect_0 (
		.ARM_A9_HPS_h2f_axi_master_awid                                        (arm_a9_hps_h2f_axi_master_awid),            //                                       ARM_A9_HPS_h2f_axi_master.awid
		.ARM_A9_HPS_h2f_axi_master_awaddr                                      (arm_a9_hps_h2f_axi_master_awaddr),          //                                                                .awaddr
		.ARM_A9_HPS_h2f_axi_master_awlen                                       (arm_a9_hps_h2f_axi_master_awlen),           //                                                                .awlen
		.ARM_A9_HPS_h2f_axi_master_awsize                                      (arm_a9_hps_h2f_axi_master_awsize),          //                                                                .awsize
		.ARM_A9_HPS_h2f_axi_master_awburst                                     (arm_a9_hps_h2f_axi_master_awburst),         //                                                                .awburst
		.ARM_A9_HPS_h2f_axi_master_awlock                                      (arm_a9_hps_h2f_axi_master_awlock),          //                                                                .awlock
		.ARM_A9_HPS_h2f_axi_master_awcache                                     (arm_a9_hps_h2f_axi_master_awcache),         //                                                                .awcache
		.ARM_A9_HPS_h2f_axi_master_awprot                                      (arm_a9_hps_h2f_axi_master_awprot),          //                                                                .awprot
		.ARM_A9_HPS_h2f_axi_master_awvalid                                     (arm_a9_hps_h2f_axi_master_awvalid),         //                                                                .awvalid
		.ARM_A9_HPS_h2f_axi_master_awready                                     (arm_a9_hps_h2f_axi_master_awready),         //                                                                .awready
		.ARM_A9_HPS_h2f_axi_master_wid                                         (arm_a9_hps_h2f_axi_master_wid),             //                                                                .wid
		.ARM_A9_HPS_h2f_axi_master_wdata                                       (arm_a9_hps_h2f_axi_master_wdata),           //                                                                .wdata
		.ARM_A9_HPS_h2f_axi_master_wstrb                                       (arm_a9_hps_h2f_axi_master_wstrb),           //                                                                .wstrb
		.ARM_A9_HPS_h2f_axi_master_wlast                                       (arm_a9_hps_h2f_axi_master_wlast),           //                                                                .wlast
		.ARM_A9_HPS_h2f_axi_master_wvalid                                      (arm_a9_hps_h2f_axi_master_wvalid),          //                                                                .wvalid
		.ARM_A9_HPS_h2f_axi_master_wready                                      (arm_a9_hps_h2f_axi_master_wready),          //                                                                .wready
		.ARM_A9_HPS_h2f_axi_master_bid                                         (arm_a9_hps_h2f_axi_master_bid),             //                                                                .bid
		.ARM_A9_HPS_h2f_axi_master_bresp                                       (arm_a9_hps_h2f_axi_master_bresp),           //                                                                .bresp
		.ARM_A9_HPS_h2f_axi_master_bvalid                                      (arm_a9_hps_h2f_axi_master_bvalid),          //                                                                .bvalid
		.ARM_A9_HPS_h2f_axi_master_bready                                      (arm_a9_hps_h2f_axi_master_bready),          //                                                                .bready
		.ARM_A9_HPS_h2f_axi_master_arid                                        (arm_a9_hps_h2f_axi_master_arid),            //                                                                .arid
		.ARM_A9_HPS_h2f_axi_master_araddr                                      (arm_a9_hps_h2f_axi_master_araddr),          //                                                                .araddr
		.ARM_A9_HPS_h2f_axi_master_arlen                                       (arm_a9_hps_h2f_axi_master_arlen),           //                                                                .arlen
		.ARM_A9_HPS_h2f_axi_master_arsize                                      (arm_a9_hps_h2f_axi_master_arsize),          //                                                                .arsize
		.ARM_A9_HPS_h2f_axi_master_arburst                                     (arm_a9_hps_h2f_axi_master_arburst),         //                                                                .arburst
		.ARM_A9_HPS_h2f_axi_master_arlock                                      (arm_a9_hps_h2f_axi_master_arlock),          //                                                                .arlock
		.ARM_A9_HPS_h2f_axi_master_arcache                                     (arm_a9_hps_h2f_axi_master_arcache),         //                                                                .arcache
		.ARM_A9_HPS_h2f_axi_master_arprot                                      (arm_a9_hps_h2f_axi_master_arprot),          //                                                                .arprot
		.ARM_A9_HPS_h2f_axi_master_arvalid                                     (arm_a9_hps_h2f_axi_master_arvalid),         //                                                                .arvalid
		.ARM_A9_HPS_h2f_axi_master_arready                                     (arm_a9_hps_h2f_axi_master_arready),         //                                                                .arready
		.ARM_A9_HPS_h2f_axi_master_rid                                         (arm_a9_hps_h2f_axi_master_rid),             //                                                                .rid
		.ARM_A9_HPS_h2f_axi_master_rdata                                       (arm_a9_hps_h2f_axi_master_rdata),           //                                                                .rdata
		.ARM_A9_HPS_h2f_axi_master_rresp                                       (arm_a9_hps_h2f_axi_master_rresp),           //                                                                .rresp
		.ARM_A9_HPS_h2f_axi_master_rlast                                       (arm_a9_hps_h2f_axi_master_rlast),           //                                                                .rlast
		.ARM_A9_HPS_h2f_axi_master_rvalid                                      (arm_a9_hps_h2f_axi_master_rvalid),          //                                                                .rvalid
		.ARM_A9_HPS_h2f_axi_master_rready                                      (arm_a9_hps_h2f_axi_master_rready),          //                                                                .rready
		.System_PLL_sys_clk_clk                                                (system_pll_sys_clk_clk),                    //                                              System_PLL_sys_clk.clk
		.ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),        // ARM_A9_HPS_h2f_axi_master_agent_clk_reset_reset_bridge_in_reset.reset
		.inst_sram_reset2_reset_bridge_in_reset_reset                          (rst_controller_001_reset_out_reset),        //                          inst_sram_reset2_reset_bridge_in_reset.reset
		.done_sram_s2_address                                                  (mm_interconnect_0_done_sram_s2_address),    //                                                    done_sram_s2.address
		.done_sram_s2_write                                                    (mm_interconnect_0_done_sram_s2_write),      //                                                                .write
		.done_sram_s2_readdata                                                 (mm_interconnect_0_done_sram_s2_readdata),   //                                                                .readdata
		.done_sram_s2_writedata                                                (mm_interconnect_0_done_sram_s2_writedata),  //                                                                .writedata
		.done_sram_s2_chipselect                                               (mm_interconnect_0_done_sram_s2_chipselect), //                                                                .chipselect
		.done_sram_s2_clken                                                    (mm_interconnect_0_done_sram_s2_clken),      //                                                                .clken
		.inst_sram_s2_address                                                  (mm_interconnect_0_inst_sram_s2_address),    //                                                    inst_sram_s2.address
		.inst_sram_s2_write                                                    (mm_interconnect_0_inst_sram_s2_write),      //                                                                .write
		.inst_sram_s2_readdata                                                 (mm_interconnect_0_inst_sram_s2_readdata),   //                                                                .readdata
		.inst_sram_s2_writedata                                                (mm_interconnect_0_inst_sram_s2_writedata),  //                                                                .writedata
		.inst_sram_s2_byteenable                                               (mm_interconnect_0_inst_sram_s2_byteenable), //                                                                .byteenable
		.inst_sram_s2_chipselect                                               (mm_interconnect_0_inst_sram_s2_chipselect), //                                                                .chipselect
		.inst_sram_s2_clken                                                    (mm_interconnect_0_inst_sram_s2_clken),      //                                                                .clken
		.sram_0_s2_address                                                     (mm_interconnect_0_sram_0_s2_address),       //                                                       sram_0_s2.address
		.sram_0_s2_write                                                       (mm_interconnect_0_sram_0_s2_write),         //                                                                .write
		.sram_0_s2_readdata                                                    (mm_interconnect_0_sram_0_s2_readdata),      //                                                                .readdata
		.sram_0_s2_writedata                                                   (mm_interconnect_0_sram_0_s2_writedata),     //                                                                .writedata
		.sram_0_s2_byteenable                                                  (mm_interconnect_0_sram_0_s2_byteenable),    //                                                                .byteenable
		.sram_0_s2_chipselect                                                  (mm_interconnect_0_sram_0_s2_chipselect),    //                                                                .chipselect
		.sram_0_s2_clken                                                       (mm_interconnect_0_sram_0_s2_clken),         //                                                                .clken
		.sram_1_s2_address                                                     (mm_interconnect_0_sram_1_s2_address),       //                                                       sram_1_s2.address
		.sram_1_s2_write                                                       (mm_interconnect_0_sram_1_s2_write),         //                                                                .write
		.sram_1_s2_readdata                                                    (mm_interconnect_0_sram_1_s2_readdata),      //                                                                .readdata
		.sram_1_s2_writedata                                                   (mm_interconnect_0_sram_1_s2_writedata),     //                                                                .writedata
		.sram_1_s2_byteenable                                                  (mm_interconnect_0_sram_1_s2_byteenable),    //                                                                .byteenable
		.sram_1_s2_chipselect                                                  (mm_interconnect_0_sram_1_s2_chipselect),    //                                                                .chipselect
		.sram_1_s2_clken                                                       (mm_interconnect_0_sram_1_s2_clken),         //                                                                .clken
		.sram_2_s2_address                                                     (mm_interconnect_0_sram_2_s2_address),       //                                                       sram_2_s2.address
		.sram_2_s2_write                                                       (mm_interconnect_0_sram_2_s2_write),         //                                                                .write
		.sram_2_s2_readdata                                                    (mm_interconnect_0_sram_2_s2_readdata),      //                                                                .readdata
		.sram_2_s2_writedata                                                   (mm_interconnect_0_sram_2_s2_writedata),     //                                                                .writedata
		.sram_2_s2_byteenable                                                  (mm_interconnect_0_sram_2_s2_byteenable),    //                                                                .byteenable
		.sram_2_s2_chipselect                                                  (mm_interconnect_0_sram_2_s2_chipselect),    //                                                                .chipselect
		.sram_2_s2_clken                                                       (mm_interconnect_0_sram_2_s2_clken),         //                                                                .clken
		.sram_3_s2_address                                                     (mm_interconnect_0_sram_3_s2_address),       //                                                       sram_3_s2.address
		.sram_3_s2_write                                                       (mm_interconnect_0_sram_3_s2_write),         //                                                                .write
		.sram_3_s2_readdata                                                    (mm_interconnect_0_sram_3_s2_readdata),      //                                                                .readdata
		.sram_3_s2_writedata                                                   (mm_interconnect_0_sram_3_s2_writedata),     //                                                                .writedata
		.sram_3_s2_byteenable                                                  (mm_interconnect_0_sram_3_s2_byteenable),    //                                                                .byteenable
		.sram_3_s2_chipselect                                                  (mm_interconnect_0_sram_3_s2_chipselect),    //                                                                .chipselect
		.sram_3_s2_clken                                                       (mm_interconnect_0_sram_3_s2_clken),         //                                                                .clken
		.sram_4_s2_address                                                     (mm_interconnect_0_sram_4_s2_address),       //                                                       sram_4_s2.address
		.sram_4_s2_write                                                       (mm_interconnect_0_sram_4_s2_write),         //                                                                .write
		.sram_4_s2_readdata                                                    (mm_interconnect_0_sram_4_s2_readdata),      //                                                                .readdata
		.sram_4_s2_writedata                                                   (mm_interconnect_0_sram_4_s2_writedata),     //                                                                .writedata
		.sram_4_s2_byteenable                                                  (mm_interconnect_0_sram_4_s2_byteenable),    //                                                                .byteenable
		.sram_4_s2_chipselect                                                  (mm_interconnect_0_sram_4_s2_chipselect),    //                                                                .chipselect
		.sram_4_s2_clken                                                       (mm_interconnect_0_sram_4_s2_clken),         //                                                                .clken
		.sram_5_s2_address                                                     (mm_interconnect_0_sram_5_s2_address),       //                                                       sram_5_s2.address
		.sram_5_s2_write                                                       (mm_interconnect_0_sram_5_s2_write),         //                                                                .write
		.sram_5_s2_readdata                                                    (mm_interconnect_0_sram_5_s2_readdata),      //                                                                .readdata
		.sram_5_s2_writedata                                                   (mm_interconnect_0_sram_5_s2_writedata),     //                                                                .writedata
		.sram_5_s2_byteenable                                                  (mm_interconnect_0_sram_5_s2_byteenable),    //                                                                .byteenable
		.sram_5_s2_chipselect                                                  (mm_interconnect_0_sram_5_s2_chipselect),    //                                                                .chipselect
		.sram_5_s2_clken                                                       (mm_interconnect_0_sram_5_s2_clken),         //                                                                .clken
		.sram_6_s2_address                                                     (mm_interconnect_0_sram_6_s2_address),       //                                                       sram_6_s2.address
		.sram_6_s2_write                                                       (mm_interconnect_0_sram_6_s2_write),         //                                                                .write
		.sram_6_s2_readdata                                                    (mm_interconnect_0_sram_6_s2_readdata),      //                                                                .readdata
		.sram_6_s2_writedata                                                   (mm_interconnect_0_sram_6_s2_writedata),     //                                                                .writedata
		.sram_6_s2_byteenable                                                  (mm_interconnect_0_sram_6_s2_byteenable),    //                                                                .byteenable
		.sram_6_s2_chipselect                                                  (mm_interconnect_0_sram_6_s2_chipselect),    //                                                                .chipselect
		.sram_6_s2_clken                                                       (mm_interconnect_0_sram_6_s2_clken),         //                                                                .clken
		.sram_7_s2_address                                                     (mm_interconnect_0_sram_7_s2_address),       //                                                       sram_7_s2.address
		.sram_7_s2_write                                                       (mm_interconnect_0_sram_7_s2_write),         //                                                                .write
		.sram_7_s2_readdata                                                    (mm_interconnect_0_sram_7_s2_readdata),      //                                                                .readdata
		.sram_7_s2_writedata                                                   (mm_interconnect_0_sram_7_s2_writedata),     //                                                                .writedata
		.sram_7_s2_byteenable                                                  (mm_interconnect_0_sram_7_s2_byteenable),    //                                                                .byteenable
		.sram_7_s2_chipselect                                                  (mm_interconnect_0_sram_7_s2_chipselect),    //                                                                .chipselect
		.sram_7_s2_clken                                                       (mm_interconnect_0_sram_7_s2_clken),         //                                                                .clken
		.sram_8_s2_address                                                     (mm_interconnect_0_sram_8_s2_address),       //                                                       sram_8_s2.address
		.sram_8_s2_write                                                       (mm_interconnect_0_sram_8_s2_write),         //                                                                .write
		.sram_8_s2_readdata                                                    (mm_interconnect_0_sram_8_s2_readdata),      //                                                                .readdata
		.sram_8_s2_writedata                                                   (mm_interconnect_0_sram_8_s2_writedata),     //                                                                .writedata
		.sram_8_s2_byteenable                                                  (mm_interconnect_0_sram_8_s2_byteenable),    //                                                                .byteenable
		.sram_8_s2_chipselect                                                  (mm_interconnect_0_sram_8_s2_chipselect),    //                                                                .chipselect
		.sram_8_s2_clken                                                       (mm_interconnect_0_sram_8_s2_clken)          //                                                                .clken
	);

	Computer_System_irq_mapper irq_mapper (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq0_irq)  //    sender.irq
	);

	Computer_System_irq_mapper irq_mapper_001 (
		.clk        (),                        //       clk.clk
		.reset      (),                        // clk_reset.reset
		.sender_irq (arm_a9_hps_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),      // reset_in1.reset
		.clk            (pll_0_outclk0_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),            // reset_in0.reset
		.reset_in1      (system_pll_reset_source_reset),          // reset_in1.reset
		.clk            (system_pll_sys_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~arm_a9_hps_h2f_reset_reset),        // reset_in0.reset
		.clk            (system_pll_sys_clk_clk),             //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
